module main

fn main() {
	// String literal printing
	println('hello')

	// String variable
	s := 'world'
	println(s)

	// String length
	println(s.len)

	// String concatenation
	greeting := 'hello' + ' ' + 'world'
	println(greeting)
	println(greeting.len)
}
