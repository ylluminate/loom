module main

fn main() {
	a := 100
	b := 7
	println(a + b)
	println(a - b)
	println(a * b)
	println(a / b)
	println(a % b)
}
