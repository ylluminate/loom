module main

fn main() {
	println(42)
}
